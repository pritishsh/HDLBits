module top_module( 
    input a, 
    input b, 
    output out );
    xnor xnor1 (out,a,b);
endmodule
