module top_module( 
    input a, 
    input b, 
    output out );
    nor nor1 (out,a,b);
endmodule
